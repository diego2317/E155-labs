// Author: Diego Weiss
// Email: dweiss@hmc.edu
// Date: 9/15/25
// This package defines statetypes to improve code readability
package state;
	// define variable type for state
	typedef enum logic [4:0] {R0, R1, R2, R3, B0, B1, B2, B3, D0, D1, D2, D3, P0, P1, P2, P3, W0, W1, W2, W3} statetype;
endpackage