// Author: Diego Weiss
// Email: dweiss@hmc.edu
// Date: 9/13/25
// This module is a top-level testbench for my implementation of E155 Lab 3
module lab3_dw_tb();


endmodule